`timescale 1ns / 1ns
`include "mux41_4.v"

module mux41_4_tb;
    wire[3:0] Y;
    reg[3:0] w0, w1, w2, w3;
    reg[1:0] S;
    // mux41_4(w0,w1,w2,w3,s,y);
    mux41_4 mux(w0,w1,w2,w3,S,Y);

    initial begin
        $dumpfile("mux41_4_tb.vcd");
        $dumpvars(0, mux41_4_tb);

        w0 = 4'b0001; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b1000;
        S = 2'b00;
        #20
        w0 = 4'b0010; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b0100;
        S = 2'b01;
        #20
        w0 = 4'b0011; w1 = 4'b1010; w2 = 4'b0011; w3 = 4'b1000;
        S = 2'b10;
        #20
        w0 = 4'b0100; w1 = 4'b0010; w2 = 4'b1100; w3 = 4'b0000;
        S = 2'b00;
        #20
        w0 = 4'b0101; w1 = 4'b0010; w2 = 4'b1000; w3 = 4'b0000;
        S = 2'b11;
        #20
        w0 = 4'b0111; w1 = 4'b0010; w2 = 4'b0010; w3 = 4'b0000;
        S = 2'b00;
        #20
        w0 = 4'b1000; w1 = 4'b0010; w2 = 4'b0100; w3 = 4'b0000;
        S = 2'b10;
        #20
        w0 = 4'b1001; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b0000;
        S = 2'b01;
        #20
        w0 = 4'b1010; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b0000;
        S = 2'b11;
        #20
        w0 = 4'b1011; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b0000;
        S = 2'b01;
        #20
        w0 = 4'b1100; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b0000;
        S = 2'b00;
        #20
        w0 = 4'b1101; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b0000;
        S = 2'b10;
        #20
        w0 = 4'b1110; w1 = 4'b0010; w2 = 4'b0000; w3 = 4'b0000;
        S = 2'b00;
        #20
        
        $display("Finish test!");
        $finish;
    end
endmodule
